class packet; endclass
