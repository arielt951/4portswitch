module switch_4port (input logic clk, input logic rst_n,
  port_if port0, port_if port1, port_if port2, port_if port3);

// Use parameters and DEFINE
// Modular design with wiring

endmodule
