    Mac OS X            	   2  >     p                                      ATTR      p   �   �                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl     4   <  com.apple.quarantine �0$i    ��)     }���Nď�֠E���                                                      q/0081;69241dd4;Chrome;6E7BD442-B988-4C59-8152-4B9FBF55CF0A 