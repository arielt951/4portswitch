class agent extends component_base; function new(string n, component_base p=null); super.new(n,p); endfunction endclass
